module top_module ( 
    input p1a, p1b, p1c, p1d,
    output reg p1y,
    input p2a, p2b, p2c, p2d,
    output reg p2y );
    
    always@(p1a,p1b,p1c,p1d)
    p1y<=~(p1a&p1b&p1c&p1d);
    always@(p2a,p2b,p2c,p2d)
    p2y<=~(p2a&p2b&p2c&p2d);

endmodule
